package pkg_definitions;
parameter NBITS = 4;
typedef enum {RESET, LOAD, UP, DOWN} counter_op_e;

endpackage
