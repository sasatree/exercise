class component_base_t;
virtual simple_if vif;

function void setup_if(virtual simple_if sif);
    vif = sif;
endfunction

endclass
