`ifndef PKG_H
`define PKG_H

`include "pkg_definitions.sv"

package pkg;
import pkg_definitions::*;

`include "simple_item.sv"
`include "test_base.sv"
`include "test1.sv"
`include "test2.sv"
`include "component_base.sv"
`include "driver.sv"
`include "run_param.sv"
`include "collector.sv"
`include "testbench.sv"

endpackage

`endif
