`ifndef PKG_H
`define PKG_H

`include "pkg_definitions.sv"

package pkg;
import uvm_pkg::*;
import pkg_definitions::*;

`include "simple_item.sv"
`include "simple_sequence_load.sv"
`include "simple_sequence_up.sv"
`include "simple_sequence_down.sv"
`include "simple_sequence_base.sv"
`include "simple_sequence1.sv"
`include "simple_sequence2.sv"
`include "simple_sequencer.sv"
`include "simple_collector.sv"
`include "simple_monitor.sv"
`include "simple_driver.sv"
`include "simple_agent.sv"
`include "simple_env.sv"
`include "simple_test_base.sv"
`include "simple_test1.sv"
`include "simple_test2.sv"
`include "simple_sequence_reset.sv"
endpackage

`endif
